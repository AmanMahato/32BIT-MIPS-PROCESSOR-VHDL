----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    15:57:43 12/04/2016 
-- Design Name: 
-- Module Name:    Instr_Mem - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL; --use CONV_INTEGER

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

 
entity InstructionMemory is
	PORT  (
			 PC: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			 instruction: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)); --31-bit output
end InstructionMemory;

architecture Behavioral of InstructionMemory is

TYPE MEMORY IS ARRAY (0 TO 127) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
CONSTANT imem: MEMORY := (   X"00000000",

"00000000000000000101000000010000",--1
"00000000000000000100000000010000",--2
"00000000000000000100100000010000",--3
"00000000000000000000100000010000",--4
"00000100000100010000000001001110",--5
"00000100000100100000000000011010",--6
"00000100000100110000000000000100",--7
"00101010001010100000000000011100",--8
"00011101000010110000000000000010",--9
"00000001011001000101100000010000",--10 
"00000001011001110001100000010000",--11 
"00010100011011010000000000000011",--12
"00011000011011100000000000011101",--13 
"00000001101011100010000000010000",--14 
"00000000100000100010100000010000",--15
"00011101001011000000000000011100",--16
"00000001100001010011000000010000",--17
"00001100101011100000000000011111",--18
"00000000000000000110100000010000",--19
"00000000000001100011100000010000",--20
"00101001101011100000000000000101",--21
"00010100111011110000000000000001",--22
"00011000111100000000000000011111",--23 
"00000001111100000011100000010000",--24
"00000101101011010000000000000001",--25 
"00110000000000000000000000010101",--26 
"00100001000001000000000000000010",--27
"00100001001001110000000000011100",--28
"00000101000010000000000000000001",--29 
"00000101001010010000000000000001",--30
"00000101010010100000000000000001",--31
"00101101000100100000000000000001",--32
"00000000000000000100000000010000",--33
"00101101001100110000000000000001",--34
"00000000000000000100100000010000",--35
"00110000000000000000000000001000",--36
"00011100000000010000000000000000",--37 
"00011100000000100000000000000001",--38
"00000000000000000001100000010000",--39
"00000100000111100000000000011010",--40 
"00000000000000000010000000010000",--41
"00000000000000000010100000010000",--42 
"00011100011111110000000000000010",--43
"00000000001111110010000000010000",--44
"00011100011111110000000000000011",--45
"00000000010111110010100000010000",--46
"00000100011000110000000000000010",--47
"00101000011111100000000000011110",--48
"00000000100001010011000000010010",--49
"00000000100001010011100000010100",--50
"00000000110001110100000000010100",--51
"00001100101001110000000000011111",--52
"00000000000000000011000000010000",--53
"00000000000010000100100000010000",--54
"00101000110001110000000000000101",--55
"00010101001010100000000000000001",--56
"00011001001010110000000000011111",--57
"00000001010010110100100000010000",--58
"00000100110001100000000000000001",--59
"00110000000000000000000000110111",--60
"00011100011111110000000000000010",--61
"00000001001111110010000000010000",--62
"00000000100001010011000000010010",--63
"00000000101001000011100000010100",--64
"00000000110001110110000000010100",--65 
"00001100100001110000000000011111",--66 
"00000000000000000011000000010000",--67
"00000000000011000110100000010000",--68
"00101000110001110000000000000101",--69
"00010101101010100000000000000001",--70
"00011001101010110000000000011111",--71
"00000001010010110110100000010000",--72
"00000100110001100000000000000001",--73
"00110000000000000000000001000101",--74
"00011100011111110000000000000011",--75
"00000001101111110010100000010000",--76 
"00000100011000110000000000000010",--77
"00110000000000000000000000110000",--78
"00100000000001000000000000100000",--79
"00100000000001010000000000100001",--80
"00011100000001000000000000100000",--81
"00011100000001010000000000100001",--82
"00000100000000110000000000011000",--83
"00101000011000000000000000011110",--84
"00011100011010000000000000000011",--85
"00000000101010000011100000010001",--86
"00001100100010010000000000011111",--87
"00000000000000000100000000010000",--88
"00000000000001110101100000010000",--89
"00101001000010010000000000000101",--90
"00011001011011000000000000000001",--91
"00010101011011010000000000011111",--92
"00000001100011010101100000010000",--93
"00000101000010000000000000000001",--94
"00110000000000000000000001011010",--95
"00000000100010110100000000010010",--96 
"00000001011001000100100000010100",--97 
"00000001000010010010100000010100",--98 
"00011100011010000000000000000010",--99
"00000000100010000011000000010001",--100
"00001100101010010000000000011111",--101
"00000000000000000100000000010000",--102
"00000000000001100101000000010000",--103
"00101001000010010000000000000101",--104 
"00011001010011000000000000000001",--105
"00010101010011010000000000011111",--106
"00000001100011010101000000010000",--107 
"00000101000010000000000000000001",--108
"00110000000000000000000001101000",--109
"00000001010001010100000000010100",--110
"00000000101010100100100000010010",--111
"00000001000010010010000000010100",--112 
"00001000011000110000000000000010",--113
"00110000000000000000000001010100",--114
"00011100011010000000000000000011",--115
"00000000101010000010100000010001",--116
"00011100011010000000000000000010",--117
"00000000100010000010000000010001",--118 
"00100000000001000000000000100010",--119
"00100000000001010000000000100011",--120

"11111100000000000000000000000000",--HALT 
 X"00000000", X"00000000",
X"00000000", X"00000000", X"00000000",X"00000000"
); 

BEGIN

instruction <= imem(CONV_INTEGER(PC(6 downto 0)));

end Behavioral;


